library verilog;
use verilog.vl_types.all;
entity TestCounter is
end TestCounter;
