library verilog;
use verilog.vl_types.all;
entity TestCntSecMinHr is
end TestCntSecMinHr;
