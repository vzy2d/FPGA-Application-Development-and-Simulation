library verilog;
use verilog.vl_types.all;
entity TestAxi4Lite is
end TestAxi4Lite;
