library verilog;
use verilog.vl_types.all;
entity CombFunctions is
end CombFunctions;
