library verilog;
use verilog.vl_types.all;
entity TestSpi is
end TestSpi;
