library verilog;
use verilog.vl_types.all;
entity TestAxi4StreamFifo is
end TestAxi4StreamFifo;
