library verilog;
use verilog.vl_types.all;
entity TestScFifo is
end TestScFifo;
