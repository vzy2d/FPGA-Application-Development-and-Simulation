library verilog;
use verilog.vl_types.all;
entity TestAxi4Stream is
end TestAxi4Stream;
