library verilog;
use verilog.vl_types.all;
entity TestMem is
end TestMem;
