library verilog;
use verilog.vl_types.all;
entity PicoMmInterconnector1to3 is
end PicoMmInterconnector1to3;
