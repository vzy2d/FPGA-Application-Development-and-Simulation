library verilog;
use verilog.vl_types.all;
entity Axi4LiteMasterEg is
    port(
        start           : in     vl_logic
    );
end Axi4LiteMasterEg;
