library verilog;
use verilog.vl_types.all;
entity TestPicoMmIf is
end TestPicoMmIf;
