library verilog;
use verilog.vl_types.all;
entity Axi4sFifo is
end Axi4sFifo;
